module FINAL(
	input CLOCK_50
);
PlatformDesigner (CLOCK_50,1'b1);
endmodule